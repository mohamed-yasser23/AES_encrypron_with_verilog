module decipherDE(clk,in,out,key);

input clk;
input [127:0] in;
input [127:0] key;
output [127:0] out;
reg [3:0] count = 4'd0;
reg [127:0] reg_in,temp;
wire [127:0] ST4,ST5,ST6,invOutSHIFT,invOutSUB;
wire [128*(10+1)-1:0] RoundKeys;

Key_Generator k(key,RoundKeys);
addRoundKey K12(in , RoundKeys[127:0] , ST4);

decryptRound DE(reg_in,RoundKeys[(((128*(10+1))-1)-128*(10-count)) -:128],ST5);

Invshiftrows invrow (reg_in,invOutSHIFT);
inverseSubBytes invsub (invOutSHIFT,invOutSUB);
addRoundKey invaddkey (invOutSUB,RoundKeys[(128*(10+1)-1) -: 128],ST6);

always @ (posedge clk) begin
$display ("ST4 = %h,ST5 = %h,ST6 = %h", ST4,ST5,ST6);
$display ("invRound = %d", count);
if(count==4'd0) begin
    reg_in<=ST4;
    temp<=ST4;
    count<=count + 4'd1;
end
else if(count<4'd10) begin
    reg_in<=ST5;
    temp<=ST5;
    count<=count + 4'd1;
end
else if(count==4'd10) begin
    reg_in<=ST5;
    temp<=ST6;
    count <= 4'd0;
end
end
assign out=temp;

endmodule